`ifndef WISHBONE_MONITOR__SV
`define WISHBONE_MONITOR__SV


class wishbone_monitor extends uvm_monitor;

//To Add
 
endclass

`endif  //WISHBONE_MONITOR__SV