`ifndef TEST_LIB__SVH
`define TEST_LIB__SVH

`include "../testcases/test_loopback.sv"
`include "../testcases/test_small_packet.sv"
`include "../testcases/test_large_packet.sv"

`endif  // TEST_LIB__SVH